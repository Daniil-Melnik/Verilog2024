module Lab3(clock, z_0, z_1, z_2);
    input wire clock; // высокочастотный тактовый сигнал
    output wire z_0, z_1, z_2; // выходы функций
    wire [3:0] x_in; // входные воздействия на дешифратор
    wire [7:0] y; // связи с выходами дешифратора
    reg [24:0] clock2; // низкочастотный тактовый сигнал

    // формирование низкочастотного таактового сигнала
    lpm_counter clk1 (
        .clock(clock),  // входной тактовый сигнал
        .cnt_en(1'b1),  // включение счетчика
        .sclr(1'b0),    // сброс счетчика (по умолчанию неактивен)
        .q(clock2)      // счётчик для низкочастотного тактового сигнала
    );
    defparam clk1.lpm_width = 25; // установка ширины счётчика q в 25
    // формирование входных воздействий на дешифратор (через переполнение)
    lpm_counter clk2 (
        .clock(clock2[24]), // низкочастотный тактовый сигнал
        .cnt_en(1'b1),      // включение счётчика
        .sclr(1'b0),        // сброс счётчика (по умолчанию неактивен)
        .q(x_in)            // тестовые воздействия (инкрементация)
    );
    defparam clk2.lpm_width = 4; // ширина второго счётчика q в 4

    lpm_decode decoder ( // библиотечный дешифратор
        .data(x_in),
        .eq(y)
    );
	 
	defparam decoder.lpm_width = 3;     // ширина входной шины 3 (x2x1x0)
	defparam decoder.lpm_decodes = 8;   // ширина выходной шины 8 (0-7)

    or or4(z_0, y[0], y[3], y[4], y[5]); // сборки по ИЛИ
    or or6(z_1, y[2], y[3], y[4], y[6]);
    or or1(z_2, y[0], y[6]); 
endmodule