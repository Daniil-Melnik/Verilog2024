//`timescale 1 ns / 1 ns
module lab3_1_tb;

  parameter delay= 0;

  // образцовые логические функции
  parameter tt4 = 8'b00111001;
  parameter tt6 = 8'b01011100;
  // parameter tt1 = 8'b01000001; // корректная функция
  parameter tt1 = 8'b11111111; //некорректная функция

  reg [3:0] x_in; // переменная для входных воздействий
  wire [7:0] y_out; // внутренняя переменная для состояния дешифратора
  wire z_0, z_1, z_2; // выходы логических функций
  reg [3:0] takt;  // перенная счётчик для перебора входных воздействий

  reg chech_point; // точка контроля функции тестером
  reg error_0, error_1, error_2; // сигналы тестера об ошибках
  wire vt_0, vt_1, vt_2; // образцовые значения функций

  lab3_1  lab3_1_inst ( // вставка основного модуля
    .x_in(x_in),
    .z_0(z_0),
    .z_1(z_1),
    .z_2(z_2)
  );

  initial
  begin // формирование тестовых последовательностей
    chech_point=0; // инициализация точки контроля
    for (takt = 0; takt <= 7; takt = takt + 1) // перебор входных воздействий
    begin #10;
      x_in=takt; // установка тестового воздействия
      chech_point= # delay 1; // установка точки контроля в 1
      #3;                     // на 3 ед. модельного времени
      chech_point=0; // сброс точки контроля
    end
  end
  assign vt_0 = tt4[x_in]; // присвоение образцовых значений функций
  assign vt_1 = tt6[x_in];
  assign vt_2 = tt1[x_in];

  always @ (posedge chech_point) // на передний фронт точки контроля
  begin // проверки тестером
    error_0 = z_0 == vt_0 ? 0:1;
    error_1 = z_1 == vt_1 ? 0:1;
    error_2 = z_2 == vt_2 ? 0:1;
  end
  
endmodule